library verilog;
use verilog.vl_types.all;
entity first_nios2_system_cpu is
    port(
        A_ci_multi_clock: out    vl_logic;
        A_ci_multi_reset: out    vl_logic;
        clk             : in     vl_logic;
        d_address       : out    vl_logic_vector(27 downto 0);
        d_byteenable    : out    vl_logic_vector(3 downto 0);
        d_irq           : in     vl_logic_vector(31 downto 0);
        d_read          : out    vl_logic;
        d_readdata      : in     vl_logic_vector(31 downto 0);
        d_waitrequest   : in     vl_logic;
        d_write         : out    vl_logic;
        d_writedata     : out    vl_logic_vector(31 downto 0);
        i_address       : out    vl_logic_vector(27 downto 0);
        i_read          : out    vl_logic;
        i_readdata      : in     vl_logic_vector(31 downto 0);
        i_readdatavalid : in     vl_logic;
        i_waitrequest   : in     vl_logic;
        jtag_debug_module_address: in     vl_logic_vector(8 downto 0);
        jtag_debug_module_begintransfer: in     vl_logic;
        jtag_debug_module_byteenable: in     vl_logic_vector(3 downto 0);
        jtag_debug_module_debugaccess: in     vl_logic;
        jtag_debug_module_debugaccess_to_roms: out    vl_logic;
        jtag_debug_module_readdata: out    vl_logic_vector(31 downto 0);
        jtag_debug_module_resetrequest: out    vl_logic;
        jtag_debug_module_select: in     vl_logic;
        jtag_debug_module_write: in     vl_logic;
        jtag_debug_module_writedata: in     vl_logic_vector(31 downto 0);
        M_ci_multi_a    : out    vl_logic_vector(4 downto 0);
        M_ci_multi_b    : out    vl_logic_vector(4 downto 0);
        M_ci_multi_c    : out    vl_logic_vector(4 downto 0);
        M_ci_multi_clk_en: out    vl_logic;
        M_ci_multi_dataa: out    vl_logic_vector(31 downto 0);
        M_ci_multi_datab: out    vl_logic_vector(31 downto 0);
        M_ci_multi_done : in     vl_logic;
        M_ci_multi_estatus: out    vl_logic;
        M_ci_multi_ipending: out    vl_logic_vector(31 downto 0);
        M_ci_multi_n    : out    vl_logic_vector(7 downto 0);
        M_ci_multi_readra: out    vl_logic;
        M_ci_multi_readrb: out    vl_logic;
        M_ci_multi_result: in     vl_logic_vector(31 downto 0);
        M_ci_multi_start: out    vl_logic;
        M_ci_multi_status: out    vl_logic;
        M_ci_multi_writerc: out    vl_logic;
        reset_n         : in     vl_logic
    );
end first_nios2_system_cpu;
